�cgame_state
Game_State
q )�q}q(X
   total_timeqK�X	   snake_wonq�X   appleqcgame_object
Game_Object
q)�q}q(X   object_sizeq	KK�q
X   objects_coordinatesq]qK�K��qaubX   levelqh)�q}q(h	KK�qh]q(K K �qKK�qK<K<�qKZKZ�qKxKx�qK�K��qK�K��qK�K҆qK�K��qMM�qM,M,�qMJMJ�qMhMh�qM�M��q M�M��q!M�M��q"M�M��q#M�M��q$MM�q%M:M:�q&K K��q'KK҆q(K<K��q)KZM�q*KxM,�q+K�MJ�q,K�Mh�q-K�M��q.K�M��q/MM��q0M,M��q1MJM��q2MhM�q3M�M:�q4K Mh�q5KM��q6K<M��q7KZM��q8KxM��q9K�M��q:K�M�q;K�M:�q<eubX   frameq=M�MX�q>X	   time_leftq?KkX	   last_moveq@KX   level_numberqAKX   scoreqBKnX   snakeqCh)�qD}qE(h	KK�qFh]qG(MJKZ�qHM,KZ�qIMKZ�qJK�KZ�qKK�KZ�qLK�KZ�qMK�KZ�qNK�K<�qOK�K�qPK�K�qQK�K�qRK�K�qSMK�qTM,K�qUMJK�qVeubX   snake_crashedqW�X   speedqXKub.